module sprite_generator
   (output logic [62:0][62:0] sprite);

    // NOTE: This was the output of a more generalized sprite_generator module, for sprites with radius 31. 
    //      We used this version to decrease resource utilization.
    assign sprite = 'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111111000000000000000000000000000011111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111111000000000000000000000001111111111111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111111110000000000000111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111110000000011111111111111111111111111111111111111111111111111111110000000111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111111111111111111110000000011111111111111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111111000000000000011111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111111111111000000000000000000011111111111111111111111111111111111111111110000000000000000000001111111111111111111111111111111111111111100000000000000000000000111111111111111111111111111111111111111000000000000000000000000011111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

endmodule: sprite_generator
