//play_tone.sv                                                                                        0000644 0010361 0077556 00000002011 12773554737 014656  0                                                                                                    ustar   dpmcdona                        dpmcdona_unix                                                                                                                                                                                                          `timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/30/2016 02:46:47 PM
// Design Name: 
// Module Name: play_tone
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module counter
  #(parameter N = 32)
   (input logic clk, en, rst,
    output logic [N-1:0] count);

   always_ff @(posedge clk) begin
      if(rst) count <= 0;
      else if(en) count <= count + 1;
   end

endmodule: counter

module play_tone(
    input logic CLK100MHZ, BTND,
    input logic [0:0] SW, 
    output logic AUD_PWM,
    output logic AUD_SD
    );
    
   logic [14:0]  wave_counter;
   logic [6:0] 	 internal_counter;
    logic [15:0] value;
   logic 	clk_out, locked, play, playing;
   logic 	en_wave_counter, en_internal_counter, rst_wave_counter, rst_internal_counter;
   
   enum 	logic {init, play_tone} cs, ns;
   
   assign play = ~BTND;
    assign AUD_SD = SW;
    
    sine_wave_lookup (wave_counter, value);
   counter #(15) c0(CLK100MHZ, en_wave_counter, rst_wave_counter, wave_counter);
   counter #(7) c1(CLK100MHZ, en_internal_counter, rst_internal_counter, internal_counter);
   

   always_comb begin
      playing = 0;
      rst_wave_counter = 0;
      rst_internal_counter = 0;
      en_wave_counter = 0;
      en_internal_counter = 0;
      case(cs)
	init: begin
	   rst_wave_counter = 1;
	   rst_internal_counter = 1;
	   AUD_PWM = 0;
	end
	play_tone: begin
	   if (wave_counter == 'd1775) playing = 0;
	   else begin
	      if (internal_counter == 7'd127) begin
		 rst_internal_counter = 1;
		 en_wave_counter = 1;
	      end
	      else begin
		 en_internal_counter = 1;
	      end
	   end
	   AUD_PWM = (value > internal_counter);
	end // case: play_tone
      endcase // case (cs)
   end // always_comb
   
   always_ff @(posedge CLK100MHZ) begin
      if (play) cs <= play_tone;
      else if (~play && ~playing) cs <= init;
   end
   /*
    always_ff @(posedge CLK100MHZ) begin
        if (wave_counter == 'd1775) begin
            wave_counter <= 'd0;
            internal_counter <= 'd0;
        end
        else begin
            if (internal_counter == 7'd127) begin
                wave_counter <= wave_counter + 11'b1;
                internal_counter <= 'd0;
            end
            else begin
                wave_counter <= wave_counter;
                internal_counter <= internal_counter + 6'b1;
            end
        end
        AUD_PWM <= (value > internal_counter);
    end
    */
endmodule: play_tone

module sine_wave_lookup (input logic [10:0] index, output logic [6:0] value);
 
logic [1775:0][6:0] vals = {7'd0,7'd0,7'd0,7'd0,7'd0,7'd1,7'd1,7'd1,7'd1,7'd2,7'd2,7'd2,7'd2,7'd2,7'd3,7'd3,7'd3,7'd3,7'd4,
7'd4,7'd4,7'd4,7'd4,7'd5,7'd5,7'd5,7'd5,7'd6,7'd6,7'd6,7'd6,7'd7,7'd7,7'd7,7'd7,7'd7,7'd8,7'd8,7'd8,7'd8,7'd9,7'd9,7'd9,
7'd9,7'd9,7'd10,7'd10,7'd10,7'd10,7'd11,7'd11,7'd11,7'd11,7'd11,7'd12,7'd12,7'd12,7'd12,7'd13,7'd13,7'd13,7'd13,7'd14,
7'd14,7'd14,7'd14,7'd14,7'd15,7'd15,7'd15,7'd15,7'd16,7'd16,7'd16,7'd16,7'd16,7'd17,7'd17,7'd17,7'd17,7'd18,7'd18,7'd18,
7'd18,7'd18,7'd19,7'd19,7'd19,7'd19,7'd20,7'd20,7'd20,7'd20,7'd20,7'd21,7'd21,7'd21,7'd21,7'd22,7'd22,7'd22,7'd22,7'd22,
7'd23,7'd23,7'd23,7'd23,7'd24,7'd24,7'd24,7'd24,7'd24,7'd25,7'd25,7'd25,7'd25,7'd26,7'd26,7'd26,7'd26,7'd26,7'd27,7'd27,
7'd27,7'd27,7'd28,7'd28,7'd28,7'd28,7'd28,7'd29,7'd29,7'd29,7'd29,7'd30,7'd30,7'd30,7'd30,7'd30,7'd31,7'd31,7'd31,7'd31,
7'd32,7'd32,7'd32,7'd32,7'd32,7'd33,7'd33,7'd33,7'd33,7'd34,7'd34,7'd34,7'd34,7'd34,7'd35,7'd35,7'd35,7'd35,7'd35,7'd36,
7'd36,7'd36,7'd36,7'd37,7'd37,7'd37,7'd37,7'd37,7'd38,7'd38,7'd38,7'd38,7'd38,7'd39,7'd39,7'd39,7'd39,7'd40,7'd40,7'd40,
7'd40,7'd40,7'd41,7'd41,7'd41,7'd41,7'd42,7'd42,7'd42,7'd42,7'd42,7'd43,7'd43,7'd43,7'd43,7'd43,7'd44,7'd44,7'd44,7'd44,
7'd44,7'd45,7'd45,7'd45,7'd45,7'd46,7'd46,7'd46,7'd46,7'd46,7'd47,7'd47,7'd47,7'd47,7'd47,7'd48,7'd48,7'd48,7'd48,7'd48,
7'd49,7'd49,7'd49,7'd49,7'd50,7'd50,7'd50,7'd50,7'd50,7'd51,7'd51,7'd51,7'd51,7'd51,7'd52,7'd52,7'd52,7'd52,7'd52,7'd53,
7'd53,7'd53,7'd53,7'd53,7'd54,7'd54,7'd54,7'd54,7'd54,7'd55,7'd55,7'd55,7'd55,7'd56,7'd56,7'd56,7'd56,7'd56,7'd57,7'd57,
7'd57,7'd57,7'd57,7'd58,7'd58,7'd58,7'd58,7'd58,7'd59,7'd59,7'd59,7'd59,7'd59,7'd60,7'd60,7'd60,7'd60,7'd60,7'd61,7'd61,
7'd61,7'd61,7'd61,7'd62,7'd62,7'd62,7'd62,7'd62,7'd63,7'd63,7'd63,7'd63,7'd63,7'd63,7'd64,7'd64,7'd64,7'd64,7'd64,7'd65,
7'd65,7'd65,7'd65,7'd65,7'd66,7'd66,7'd66,7'd66,7'd66,7'd67,7'd67,7'd67,7'd67,7'd67,7'd68,7'd68,7'd68,7'd68,7'd68,7'd69,
7'd69,7'd69,7'd69,7'd69,7'd69,7'd70,7'd70,7'd70,7'd70,7'd70,7'd71,7'd71,7'd71,7'd71,7'd71,7'd72,7'd72,7'd72,7'd72,7'd72,
7'd72,7'd73,7'd73,7'd73,7'd73,7'd73,7'd74,7'd74,7'd74,7'd74,7'd74,7'd75,7'd75,7'd75,7'd75,7'd75,7'd75,7'd76,7'd76,7'd76,
7'd76,7'd76,7'd77,7'd77,7'd77,7'd77,7'd77,7'd77,7'd78,7'd78,7'd78,7'd78,7'd78,7'd78,7'd79,7'd79,7'd79,7'd79,7'd79,7'd80,
7'd80,7'd80,7'd80,7'd80,7'd80,7'd81,7'd81,7'd81,7'd81,7'd81,7'd81,7'd82,7'd82,7'd82,7'd82,7'd82,7'd83,7'd83,7'd83,7'd83,
7'd83,7'd83,7'd84,7'd84,7'd84,7'd84,7'd84,7'd84,7'd85,7'd85,7'd85,7'd85,7'd85,7'd85,7'd86,7'd86,7'd86,7'd86,7'd86,7'd86,
7'd87,7'd87,7'd87,7'd87,7'd87,7'd87,7'd88,7'd88,7'd88,7'd88,7'd88,7'd88,7'd89,7'd89,7'd89,7'd89,7'd89,7'd89,7'd90,7'd90,
7'd90,7'd90,7'd90,7'd90,7'd90,7'd91,7'd91,7'd91,7'd91,7'd91,7'd91,7'd92,7'd92,7'd92,7'd92,7'd92,7'd92,7'd93,7'd93,7'd93,
7'd93,7'd93,7'd93,7'd93,7'd94,7'd94,7'd94,7'd94,7'd94,7'd94,7'd95,7'd95,7'd95,7'd95,7'd95,7'd95,7'd95,7'd96,7'd96,7'd96,
7'd96,7'd96,7'd96,7'd96,7'd97,7'd97,7'd97,7'd97,7'd97,7'd97,7'd98,7'd98,7'd98,7'd98,7'd98,7'd98,7'd98,7'd99,7'd99,7'd99,
7'd99,7'd99,7'd99,7'd99,7'd100,7'd100,7'd100,7'd100,7'd100,7'd100,7'd100,7'd100,7'd101,7'd101,7'd101,7'd101,7'd101,7'd101,
7'd101,7'd102,7'd102,7'd102,7'd102,7'd102,7'd102,7'd102,7'd103,7'd103,7'd103,7'd103,7'd103,7'd103,7'd103,7'd103,7'd104,
7'd104,7'd104,7'd104,7'd104,7'd104,7'd104,7'd105,7'd105,7'd105,7'd105,7'd105,7'd105,7'd105,7'd105,7'd106,7'd106,7'd106,
7'd106,7'd106,7'd106,7'd106,7'd106,7'd107,7'd107,7'd107,7'd107,7'd107,7'd107,7'd107,7'd107,7'd108,7'd108,7'd108,7'd108,
7'd108,7'd108,7'd108,7'd108,7'd108,7'd109,7'd109,7'd109,7'd109,7'd109,7'd109,7'd109,7'd109,7'd110,7'd110,7'd110,7'd110,
7'd110,7'd110,7'd110,7'd110,7'd110,7'd111,7'd111,7'd111,7'd111,7'd111,7'd111,7'd111,7'd111,7'd111,7'd112,7'd112,7'd112,7'd112,7'd112,7'd112,7'd112,7'd112,7'd112,7'd113,7'd113,7'd113,7'd113,7'd113,7'd113,7'd113,7'd113,7'd113,7'd113,7'd114,7'd114,7'd114,7'd114,7'd114,7'd114,7'd114,7'd114,7'd114,7'd114,7'd115,7'd115,7'd115,7'd115,7'd115,7'd115,7'd115,7'd115,7'd115,7'd115,7'd116,7'd116,7'd116,7'd116,7'd116,7'd116,7'd116,7'd116,7'd116,7'd116,7'd117,7'd117,7'd117,7'd117,7'd117,7'd117,7'd117,7'd117,7'd117,7'd117,7'd117,7'd117,7'd118,7'd118,7'd118,7'd118,7'd118,7'd118,7'd118,7'd118,7'd118,7'd118,7'd118,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd128,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd127,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd126,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd125,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd124,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd123,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd122,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd121,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd120,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd119,7'd118,7'd118,7'd118,7'd118,7'd118,7'd118,7'd118,7'd118,7'd118,7'd118,7'd118,7'd117,7'd117,7'd117,7'd117,7'd117,7'd117,7'd117,7'd117,7'd117,7'd117,7'd117,7'd117,7'd116,7'd116,7'd116,7'd116,7'd116,7'd116,7'd116,7'd116,7'd116,7'd116,7'd115,7'd115,7'd115,7'd115,7'd115,7'd115,7'd115,7'd115,7'd115,7'd115,7'd114,7'd114,7'd114,7'd114,7'd114,7'd114,7'd114,7'd114,7'd114,7'd114,7'd113,7'd113,7'd113,7'd113,7'd113,7'd113,7'd113,7'd113,7'd113,7'd113,7'd112,7'd112,7'd112,7'd112,7'd112,7'd112,7'd112,7'd112,7'd112,7'd111,7'd111,7'd111,7'd111,7'd111,7'd111,7'd111,7'd111,7'd111,7'd110,7'd110,7'd110,7'd110,7'd110,7'd110,7'd110,7'd110,7'd110,7'd109,7'd109,7'd109,7'd109,7'd109,7'd109,7'd109,7'd109,7'd108,7'd108,7'd108,7'd108,7'd108,7'd108,7'd108,7'd108,7'd108,7'd107,7'd107,7'd107,7'd107,7'd107,7'd107,7'd107,7'd107,7'd106,7'd106,7'd106,7'd106,7'd106,7'd106,7'd106,7'd106,7'd105,7'd105,7'd105,7'd105,7'd105,7'd105,7'd105,7'd105,7'd104,7'd104,7'd104,7'd104,7'd104,7'd104,7'd104,7'd103,7'd103,7'd103,7'd103,7'd103,7'd103,7'd103,7'd103,7'd102,7'd102,7'd102,7'd102,7'd102,7'd102,7'd102,7'd101,7'd101,7'd101,7'd101,7'd101,7'd101,7'd101,7'd100,7'd100,7'd100,7'd100,7'd100,7'd100,7'd100,7'd100,7'd99,7'd99,7'd99,7'd99,7'd99,7'd99,7'd99,7'd98,7'd98,7'd98,7'd98,7'd98,7'd98,7'd98,7'd97,7'd97,7'd97,7'd97,7'd97,7'd97,7'd96,7'd96,7'd96,7'd96,7'd96,7'd96,7'd96,7'd95,7'd95,7'd95,7'd95,7'd95,7'd95,7'd95,7'd94,7'd94,7'd94,7'd94,7'd94,7'd94,7'd93,7'd93,7'd93,7'd93,7'd93,7'd93,7'd93,7'd92,7'd92,7'd92,7'd92,7'd92,7'd92,7'd91,7'd91,7'd91,7'd91,7'd91,7'd91,7'd90,7'd90,7'd90,7'd90,7'd90,7'd90,7'd90,7'd89,7'd89,7'd89,7'd89,7'd89,7'd89,7'd88,7'd88,7'd88,7'd88,7'd88,7'd88,7'd87,7'd87,7'd87,7'd87,7'd87,7'd87,7'd86,7'd86,7'd86,7'd86,7'd86,7'd86,7'd85,7'd85,7'd85,7'd85,7'd85,7'd85,7'd84,7'd84,7'd84,7'd84,7'd84,7'd84,7'd83,7'd83,7'd83,7'd83,7'd83,7'd83,7'd82,7'd82,7'd82,7'd82,7'd82,7'd81,7'd81,7'd81,7'd81,7'd81,7'd81,7'd80,7'd80,7'd80,7'd80,7'd80,7'd80,7'd79,7'd79,7'd79,7'd79,7'd79,7'd78,7'd78,7'd78,7'd78,7'd78,7'd78,7'd77,7'd77,7'd77,7'd77,7'd77,7'd77,7'd76,7'd76,7'd76,7'd76,7'd76,7'd75,7'd75,7'd75,7'd75,7'd75,7'd75,7'd74,7'd74,7'd74,7'd74,7'd74,7'd73,7'd73,7'd73,7'd73,7'd73,7'd72,7'd72,7'd72,7'd72,7'd72,7'd72,7'd71,7'd71,7'd71,7'd71,7'd71,7'd70,7'd70,7'd70,7'd70,7'd70,7'd69,7'd69,7'd69,7'd69,7'd69,7'd69,7'd68,7'd68,7'd68,7'd68,7'd68,7'd67,7'd67,7'd67,7'd67,7'd67,7'd66,7'd66,7'd66,7'd66,7'd66,7'd65,7'd65,7'd65,7'd65,7'd65,7'd64,7'd64,7'd64,7'd64,7'd64,7'd64,7'd63,7'd63,7'd63,7'd63,7'd63,7'd62,7'd62,7'd62,7'd62,7'd62,7'd61,7'd61,7'd61,7'd61,7'd61,7'd60,7'd60,7'd60,7'd60,7'd60,7'd59,7'd59,7'd59,7'd59,7'd59,7'd58,7'd58,7'd58,7'd58,7'd58,7'd57,7'd57,7'd57,7'd57,7'd57,7'd56,7'd56,7'd56,7'd56,7'd56,7'd55,7'd55,7'd55,7'd55,7'd54,7'd54,7'd54,7'd54,7'd54,7'd53,7'd53,7'd53,7'd53,7'd53,7'd52,7'd52,7'd52,7'd52,7'd52,7'd51,7'd51,7'd51,7'd51,7'd51,7'd50,7'd50,7'd50,7'd50,7'd50,7'd49,7'd49,7'd49,7'd49,7'd48,7'd48,7'd48,7'd48,7'd48,7'd47,7'd47,7'd47,7'd47,7'd47,7'd46,7'd46,7'd46,7'd46,7'd46,7'd45,7'd45,7'd45,7'd45,7'd44,7'd44,7'd44,7'd44,7'd44,7'd43,7'd43,7'd43,7'd43,7'd43,7'd42,7'd42,7'd42,7'd42,7'd42,7'd41,7'd41,7'd41,7'd41,7'd40,7'd40,7'd40,7'd40,7'd40,7'd39,7'd39,7'd39,7'd39,7'd38,7'd38,7'd38,7'd38,7'd38,7'd37,7'd37,7'd37,7'd37,7'd37,7'd36,7'd36,7'd36,7'd36,7'd35,7'd35,7'd35,7'd35,7'd35,7'd34,7'd34,7'd34,7'd34,7'd34,7'd33,7'd33,7'd33,7'd33,7'd32,7'd32,7'd32,7'd32,7'd32,7'd31,7'd31,7'd31,7'd31,7'd30,7'd30,7'd30,7'd30,7'd30,7'd29,7'd29,7'd29,7'd29,7'd28,7'd28,7'd28,7'd28,7'd28,7'd27,7'd27,7'd27,7'd27,7'd26,7'd26,7'd26,7'd26,7'd26,7'd25,7'd25,7'd25,7'd25,7'd24,7'd24,7'd24,7'd24,7'd24,7'd23,7'd23,7'd23,7'd23,7'd22,7'd22,7'd22,7'd22,7'd22,7'd21,7'd21,7'd21,7'd21,7'd20,7'd20,7'd20,7'd20,7'd20,7'd19,7'd19,7'd19,7'd19,7'd18,7'd18,7'd18,7'd18,7'd18,7'd17,7'd17,7'd17,7'd17,7'd16,7'd16,7'd16,7'd16,7'd16,7'd15,7'd15,7'd15,7'd15,7'd14,7'd14,7'd14,7'd14,7'd14,7'd13,7'd13,7'd13,7'd13,7'd12,7'd12,7'd12,7'd12,7'd11,7'd11,7'd11,7'd11,7'd11,7'd10,7'd10,7'd10,7'd10,7'd9,7'd9,7'd9,7'd9,7'd9,7'd8,7'd8,7'd8,7'd8,7'd7,7'd7,7'd7,7'd7,7'd7,7'd6,7'd6,7'd6,7'd6,7'd5,7'd5,7'd5,7'd5,7'd4,7'd4,7'd4,7'd4,7'd4,7'd3,7'd3,7'd3,7'd3,7'd2,7'd2,7'd2,7'd2,7'd2,7'd1,7'd1,7'd1,7'd1,7'd0,7'd0,7'd0,7'd0};

assign value = vals[index];

endmodule: sine_wave_lookup

