`define ADD 'b00
`define SUB 'b01
`define MUL 'b10
`define DIV 'b11
